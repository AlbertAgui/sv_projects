package size_fields_package;

///////////////////
//Size parameters
parameter ADDR_WIDTH=3, OPCODE_WIDTH=1, WORD_WIDTH=8;

endpackage;
