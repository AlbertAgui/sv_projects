`ifndef TEST_SVH
`define TEST_SVH

`include "uvc/package/top_uvm_pkg/top_uvm_pkg.sv"
`include "uvc/uvm_seq/seq/seq.svh"
`include "uvc/uvm_env/env/env.svh"

`include "uvc/uvm_test/test/test.sv"

`endif