`ifndef SEQ_ITEM_SVH
`define SEQ_ITEM_SVH

`include "uvc/uvm_transaction/seq_item/seq_item.sv"

`endif