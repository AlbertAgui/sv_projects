//localparam X = 3;

package visible_pkg;

class class_a;

    logic [2:0] a;

endclass //className

endpackage