`ifndef TESTBENCH_SVH
`define TESTBENCH_SVH

`include "uvc/interface/req_resp/req_resp_if.svh"
`include "uvc/package/top_uvm_pkg/top_uvm_pkg.sv"
`include "uvc/interface/int/interface.svh"

`include "uvc/testbench/tb/testbench.sv"

`endif