module Top_soc(
  input logic a_i
);

  logic temp;

  assign temp = a_i;
  
endmodule