`ifndef UVM_TEST_PKG_SV
`define UVM_TEST_PKG_SV

package uvm_test_pkg;
	import uvm_pkg::*;
	`include "uvm_macros.svh"

	`include "ka_mem_model.sv"
	`include "seq_item.sv"
	`include "driver.sv"
	`include "sequencer.sv"
	`include "seq.sv"
	`include "agent.sv"
	`include "env.sv"
	`include "v1_test.sv"
endpackage : uvm_test_pkg

`endif