`ifndef UTILS_PKG_SV
`define UTILS_PKG_SV

package utils_pkg;
	`include "transaction_cnt_wrapper.sv"
endpackage : utils_pkg

`endif