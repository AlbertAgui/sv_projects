
parameter WORD_WIDTH=4;
parameter INDEX_WIDTH=4;
parameter OPCODE_MEM_WIDTH=1;