package alu_pkg;




endpackage
