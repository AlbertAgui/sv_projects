`ifndef DUT_TOP_SVH
`define DUT_TOP_SVH

`include "rtl/dut/queue.sv"
`include "rtl/dut/dut_top.sv"

`endif