module mod1 (
    ports
);
    
endmodule