`ifndef TOP_UVM_PKG_SV
`define TOP_UVM_PKG_SV

package top_uvm_pkg;

localparam int DATA_SIZE = 16;
localparam string CNFG = "VALID_READY";
localparam int COUNT = 6;
localparam int DEPTH = 10;

localparam int SEQ_NUM = 7;

endpackage

`endif