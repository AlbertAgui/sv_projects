`ifndef UVM_SVH
`define UVM_SVH

`include "uvc/testbench/tb/testbench.svh"
`include "uvc/uvm_test/test/test.svh"

`endif