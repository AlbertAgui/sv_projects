package wb_pkg;
  typedef struct packed {
    
  } wb_req_;
endpackage