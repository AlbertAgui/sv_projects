`ifndef TEST_SVH
`define TEST_SVH

`include "uvc/uvm_seq/seq/seq.svh"
`include "uvc/uvm_env/env/env.svh"

`include "uvc/uvm_test/test/test.sv"

`endif