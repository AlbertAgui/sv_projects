`ifndef KA_SEQ_SVH
`define KA_SEQ_SVH

`include "uvc/uvm_transaction/seq_item/seq_item.svh"

`include "uvc/uvm_seq/seq/seq.sv"

`endif