class transaction_cnt_wrapper;

	int cnt;

	function new();
		this.cnt = 0;
	endfunction : new
		
endclass : transaction_cnt_wrapper