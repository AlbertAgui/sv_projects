`ifndef ENV_SVH
`define ENV_SVH

`include "uvc/interface/int/interface.svh"
`include "uvc/uvm_agent/agent/agent.svh"

`include "uvc/uvm_env/env/env.sv"

`endif