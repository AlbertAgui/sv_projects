`ifndef AGENT_SVH
`define AGENT_SVH

`include "uvc/uvm_transaction/seq_item/seq_item.svh"
`include "uvc/uvm_sequencer/sequencer/sequencer.svh"

`include "uvc/uvm_agent/agent/driver.sv"

`include "uvc/uvm_agent/agent/agent.sv"

`endif