`ifndef KA_SEQUENCER_SVH
`define KA_SEQUENCER_SVH

`include "uvc/uvm_transaction/seq_item/seq_item.svh"

`include "uvc/uvm_sequencer/sequencer/sequencer.sv"

`endif