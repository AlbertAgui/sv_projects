`ifndef TESTBENCH_SVH
`define TESTBENCH_SVH


`include "uvc/interface/int/interface.svh"

`include "uvc/testbench/tb/testbench.sv"

`endif