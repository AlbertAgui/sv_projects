`ifndef DUT_TOP_TB_SVH
`define DUT_TOP_TB_SVH

`include "uvc/interface/int/interface.svh"
`include "rtl/dut/unit_test/dut_top_tb.sv"

`endif