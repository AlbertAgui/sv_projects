`ifndef INTERFACE_SVH
`define INTERFACE_SVH

`include "uvc/interface/int/interface.sv"

`endif