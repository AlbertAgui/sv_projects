`ifndef REQ_RESP_IF_SVH
`define REQ_RESP_IF_SVH

`include "uvc/interface/req_resp/req_resp_if.sv"

`endif