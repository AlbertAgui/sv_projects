//`include "interface.sv"

module Top_soc(
  input logic a_i
);

  /*interfacename it();
  struct_name s;

  initial begin
    taskName();
  end

  //`include "interface.sv"

  logic temp;

  always_comb begin : blockName
    it.a = 1'b1;
    $display("it.a: %d", it.a);
  end

  assign temp = a_i;*/
  
endmodule